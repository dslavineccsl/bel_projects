
module issp_64i_64o (
	source,
	probe,
	source_clk);	

	output	[63:0]	source;
	input	[63:0]	probe;
	input		source_clk;
endmodule
